module and_comb(A, B, Y);
input wire A, B;
output wire Y;

assign Y = A & B;

endmodule

module AND2(A, B, X);

input A, B;
output X;

wire real A, B, X;

assign X = A + B;

endmodule
